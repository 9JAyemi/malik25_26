
module mux_stall (
	cw_from_cu, 
	mux_op, 
	cw_from_mux);
   input [22:0] cw_from_cu;
   input mux_op;
   output [22:0] cw_from_mux;

   // Internal wires
   wire n2;

   // Generate n2
   assign n2 = mux_op; // fixed the polarity

   // Implement the multiplexing logic
   assign cw_from_mux[0] = cw_from_cu[0] & n2;
   assign cw_from_mux[1] = cw_from_cu[1] & n2;
   assign cw_from_mux[2] = cw_from_cu[2] & n2;
   assign cw_from_mux[3] = cw_from_cu[3] & n2;
   assign cw_from_mux[4] = cw_from_cu[4] & n2;
   assign cw_from_mux[5] = cw_from_cu[5] & n2;
   assign cw_from_mux[6] = cw_from_cu[6] & n2;
   assign cw_from_mux[7] = cw_from_cu[7] & n2;
   assign cw_from_mux[8] = cw_from_cu[8] & n2;
   assign cw_from_mux[9] = cw_from_cu[9] & n2;
   assign cw_from_mux[10] = cw_from_cu[10] & n2;
   assign cw_from_mux[11] = cw_from_cu[11] & n2;
   assign cw_from_mux[12] = cw_from_cu[12] & n2;
   assign cw_from_mux[13] = cw_from_cu[13] & n2;
   assign cw_from_mux[14] = cw_from_cu[14] & n2;
   assign cw_from_mux[15] = cw_from_cu[15] & n2;
   assign cw_from_mux[16] = cw_from_cu[16] & n2;
   assign cw_from_mux[17] = cw_from_cu[17] & n2;
   assign cw_from_mux[18] = cw_from_cu[18] & n2;
   assign cw_from_mux[19] = cw_from_cu[19] & n2;
   assign cw_from_mux[20] = cw_from_cu[20] & n2;
   assign cw_from_mux[21] = cw_from_cu[21] & n2;
   assign cw_from_mux[22] = cw_from_cu[22] & n2;

   // Select between the two inputs based on the mux_op value
   assign cw_from_mux = cw_from_mux; // fixed the extra mux_op in the assignment
endmodule