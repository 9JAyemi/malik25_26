module up_down_counter (
    input clk,
    input rst,
    input load,
    input up_down,
    input [2:0] data_in,
    output reg [2:0] count
);

    always @(posedge clk) begin
        if (rst) begin
            count <= 3'b0;
        end else if (load) begin
            count <= data_in;
        end else if (up_down) begin
            count <= count + 1;
        end else begin
            count <= count - 1;
        end
    end

endmodule