module byte_reversal (
    input [31:0] in,
    output reg [31:0] out
);

always @(*) begin
    out[7:0] = in[31:24];
    out[15:8] = in[23:16];
    out[23:16] = in[15:8];
    out[31:24] = in[7:0];
end

endmodule

module priority_encoder (
    input [31:0] in,
    output reg [4:0] pos // Position of the first high bit in the input
);

always @(*) begin
    case(in)
        32'b00000000000000000000000000000000: pos = 5'b00000;
        32'b00000000000000000000000000000001: pos = 5'b00001;
        32'b00000000000000000000000000000011: pos = 5'b00010;
        32'b00000000000000000000000000000111: pos = 5'b00011;
        32'b00000000000000000000000000001111: pos = 5'b00100;
        32'b00000000000000000000000000011111: pos = 5'b00101;
        32'b00000000000000000000000000111111: pos = 5'b00110;
        32'b00000000000000000000000001111111: pos = 5'b00111;
        32'b00000000000000000000000011111111: pos = 5'b01000;
        32'b00000000000000000000000111111111: pos = 5'b01001;
        32'b00000000000000000000001111111111: pos = 5'b01010;
        32'b00000000000000000000011111111111: pos = 5'b01011;
        default: pos = 5'b01111;
    endcase
end

endmodule