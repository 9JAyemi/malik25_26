module binary_counter(
    input clk,
    input rst,
    output reg [3:0] count,
    output reg max_count_reached
);

always @(posedge clk) begin
    if (rst) begin
        count <= 4'b0000;
        max_count_reached <= 1'b0;
    end else if (count == 4'b1111) begin
        count <= 4'b0000;
        max_count_reached <= 1'b1;
    end else begin
        count <= count + 1;
        max_count_reached <= 1'b0;
    end
end

endmodule