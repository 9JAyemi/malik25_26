
module v053dc2 #(
 parameter v71e305 = 0
) (
 input vf54559,
 input va4102a,
 output ve8318d
);
 assign ve8318d = vf54559 & va4102a;
endmodule
module vd0c4e5 (
 input v030ad0,
 input v27dec4,
 input v2d3366,
 output vb192d0
);
 assign vb192d0 = v27dec4 ? v030ad0 : v2d3366;
endmodule
module vfebcfe (
 input v9fb85f,
 output v9fb85f_out
);
 assign v9fb85f_out = v9fb85f;
endmodule
module vd30ca9 (
 input v9fb85f,
 output v9fb85f_out
);
 assign v9fb85f_out = ~v9fb85f;
endmodule
module v144728 #(
 parameter v573b2a = 0
) (
 input v6dda25,
 input v27dec4,
 input v92a149,
 output v4642b6
);
 localparam p0 = v573b2a;
 wire w1;
 wire w3;
 wire w6;
 wire w7;
 assign w1 = v6dda25;
 v053dc2 #(
  .v71e305(p0)
 ) v24b497 (
  .vf54559(w1),
  .va4102a(w1),
  .ve8318d(w6)
 );
 vd0c4e5 vda4b54 (
  .v030ad0(w1),
  .v27dec4(v27dec4),
  .vb192d0(w3),
  .v2d3366(v27dec4)
 );
 vfebcfe v2141a0 (
  .v9fb85f(w3)
 );
 vd0c4e5 v75d8ff (
  .v030ad0(w3),
  .v27dec4(v92a149),
  .vb192d0(w7),
  .v2d3366(v92a149)
 );
 vd30ca9 va595cf (
  .v9fb85f(w7)
 );
 assign v4642b6 = w7;
endmodule