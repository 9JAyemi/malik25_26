module decoder (
    input [2:0] in,
    output [7:0] out
);
    
    assign out = {(~in[2] & ~in[1] & ~in[0]), (~in[2] & ~in[1] & in[0]), (~in[2] & in[1] & ~in[0]), (~in[2] & in[1] & in[0]), (in[2] & ~in[1] & ~in[0]), (in[2] & ~in[1] & in[0]), (in[2] & in[1] & ~in[0]), (in[2] & in[1] & in[0])};

endmodule