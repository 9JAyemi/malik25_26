module glitch_filter (
  input in,
  input clk,
  output reg out
);

parameter n = 10; // number of clock cycles to wait
parameter t = 5; // threshold value for glitch detection
parameter v = 0; // value to output when a glitch is detected

reg [n-1:0] timer;
reg glitch_detected;
reg [1:0] input_history;
wire input_above_threshold;

assign input_above_threshold = (in > t);

always @(posedge clk) begin
  if (timer == n-1) begin
    if (glitch_detected) begin
      out <= v;
    end else begin
      out <= in;
    end
    timer <= 0;
    glitch_detected <= 0;
  end else begin
    timer <= timer + 1;
    if (input_above_threshold) begin
      input_history <= {input_history[0], 1'b1};
    end else begin
      input_history <= {input_history[0], 1'b0};
    end
    if (input_history == 2'b10) begin
      glitch_detected <= 1;
    end
  end
end

endmodule