module shift_register (
  input clk,
  input reset,
  input clear,
  input [7:0] data_in,
  output [7:0] data_out
);

  reg [7:0] shift_reg;

  always @(posedge clk) begin
    if (reset) begin
      shift_reg <= 8'b0;
    end else if (clear) begin
      shift_reg <= 8'b11111111;
    end else begin
      shift_reg <= {shift_reg[6:0], data_in};
    end
  end
  
  assign data_out = shift_reg;

endmodule
