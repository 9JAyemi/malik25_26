module sumwrap_uint16_to1_1(input CLK, input CE, input [31:0] process_input, output [15:0] process_output);
parameter INSTANCE_NAME="INST";

  wire [15:0] least_sig_bits;
  assign least_sig_bits = process_input[15:0]; // Extract the least significant 16 bits of process_input
  
  wire [15:0] most_sig_bits;
  assign most_sig_bits = process_input[31:16]; // Extract the most significant 16 bits of process_input
  
  assign process_output = ((least_sig_bits == 16'd1) ? 16'd0 : (least_sig_bits + most_sig_bits)); // If least_sig_bits == 1, output 0, else output sum of least_sig_bits and most_sig_bits
  
endmodule