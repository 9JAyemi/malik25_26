
module pipelined_JC_counter(
  input                clk,
  input                rst_n,
  output reg  [15:0]   Q
);

reg [15:0] Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9, Q10, Q11, Q12, Q13, Q14, Q15, Q16;

always @(posedge clk or negedge rst_n) begin
  if(!rst_n) begin
    Q1 <= 16'b0000000000000000;
    Q2 <= 16'b0000000000000000;
    Q3 <= 16'b0000000000000000;
    Q4 <= 16'b0000000000000000;
    Q5 <= 16'b0000000000000000;
    Q6 <= 16'b0000000000000000;
    Q7 <= 16'b0000000000000000;
    Q8 <= 16'b0000000000000000;
    Q9 <= 16'b0000000000000000;
    Q10 <= 16'b0000000000000000;
    Q11 <= 16'b0000000000000000;
    Q12 <= 16'b0000000000000000;
    Q13 <= 16'b0000000000000000;
    Q14 <= 16'b0000000000000000;
    Q15 <= 16'b0000000000000000;
    Q16 <= 16'b0000000000000000;
  end else begin
    Q1 <= Q16 ^ 1'b1;
    Q2 <= Q1 ^ 1'b1;
    Q3 <= Q2 ^ 1'b1;
    Q4 <= Q3 ^ 1'b1;
    Q5 <= Q4 ^ 1'b1;
    Q6 <= Q5 ^ 1'b1;
    Q7 <= Q6 ^ 1'b1;
    Q8 <= Q7 ^ 1'b1;
    Q9 <= Q8 ^ 1'b1;
    Q10 <= Q9 ^ 1'b1;
    Q11 <= Q10 ^ 1'b1;
    Q12 <= Q11 ^ 1'b1;
    Q13 <= Q12 ^ 1'b1;
    Q14 <= Q13 ^ 1'b1;
    Q15 <= Q14 ^ 1'b1;
    Q16 <= Q15 ^ 1'b1;

    Q <= Q16;
  end
end

endmodule
