module up_counter(clk, rst, count);
  input clk;
  input rst;
  output reg [3:0] count;

  always @(posedge clk or negedge rst) begin
    if(!rst) begin
      count <= 4'b0;
    end else begin
      count <= count + 1;
    end
  end
endmodule