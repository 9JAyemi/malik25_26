module binary_counter(
  input clk,
  input rst,
  output reg [3:0] count_out,
  output reg overflow
);

  always @(posedge clk) begin
    if (rst) begin
      count_out <= 4'b0;
      overflow <= 1'b0;
    end else if (count_out == 4'b1111) begin
      count_out <= 4'b0;
      overflow <= 1'b1;
    end else begin
      count_out <= count_out + 1;
      overflow <= 1'b0;
    end
  end

endmodule