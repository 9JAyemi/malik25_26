module xor_gate(input a, b, output out_assign);
    assign out_assign = a ^ b;
endmodule