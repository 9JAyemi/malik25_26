module hamming_code #(
  parameter n = 4, // length of data_in vector
  parameter m = 7 // length of encoded_data vector (n + log2(n) + 1)
)(
  input [n-1:0] data_in,
  output [m-1:0] encoded_data,
  output [n-1:0] corrected_data
);


// Encoding
wire [m-1:0] encoded_data_temp;
assign encoded_data_temp[0] = data_in[0] ^ data_in[1] ^ data_in[3];
assign encoded_data_temp[1] = data_in[0] ^ data_in[2] ^ data_in[3];
assign encoded_data_temp[2] = data_in[0];
assign encoded_data_temp[3] = data_in[1] ^ data_in[2] ^ data_in[3];
assign encoded_data_temp[4] = data_in[1];
assign encoded_data_temp[5] = data_in[2];
assign encoded_data_temp[6] = data_in[3];
assign encoded_data = encoded_data_temp;

// Decoding
wire [m-1:0] decoded_data_temp;
wire error;
wire [2:0] error_position;
assign error = encoded_data_temp[0] ^ encoded_data_temp[1] ^ encoded_data_temp[3] ^ encoded_data_temp[4] ^ encoded_data_temp[5] ^ encoded_data_temp[6];
assign error_position = {encoded_data_temp[0] ^ encoded_data_temp[2] ^ encoded_data_temp[4] ^ encoded_data_temp[6], encoded_data_temp[1] ^ encoded_data_temp[2] ^ encoded_data_temp[5] ^ encoded_data_temp[6], encoded_data_temp[3] ^ encoded_data_temp[4] ^ encoded_data_temp[5] ^ encoded_data_temp[6]};
assign decoded_data_temp[0] = error ? (encoded_data_temp[2] ^ (error_position == 3'b001)) : encoded_data_temp[2];
assign decoded_data_temp[1] = error ? (encoded_data_temp[4] ^ (error_position == 3'b010)) : encoded_data_temp[4];
assign decoded_data_temp[2] = error ? (encoded_data_temp[5] ^ (error_position == 3'b011)) : encoded_data_temp[5];
assign decoded_data_temp[3] = error ? (encoded_data_temp[6] ^ (error_position == 3'b100)) : encoded_data_temp[6];
assign corrected_data = decoded_data_temp;

endmodule