

module RCB_FRL_CRC_gen ( D, NewCRC);

	input [47:0] D;
	output [7:0] NewCRC;
	
	
	assign NewCRC[0] = D[46] ^ D[42] ^ D[41] ^ D[37] ^ D[36] ^ D[35] ^ D[34] ^ 
                D[33] ^ D[31] ^ D[30] ^ D[29] ^ D[27] ^ D[26] ^ D[24] ^ 
                D[20] ^ D[18] ^ D[17] ^ D[16] ^ D[15] ^ D[14] ^ D[13] ^ 
                D[8] ^ D[7] ^ D[6] ^ D[3] ^ D[1] ^ D[0];
    assign NewCRC[1] = D[47] ^ D[43] ^ D[42] ^ D[38] ^ D[37] ^ D[36] ^ D[35] ^ 
                D[34] ^ D[32] ^ D[31] ^ D[30] ^ D[28] ^ D[27] ^ D[25] ^ 
                D[21] ^ D[19] ^ D[18] ^ D[17] ^ D[16] ^ D[15] ^ D[14] ^ 
                D[9] ^ D[8] ^ D[7] ^ D[4] ^ D[2] ^ D[1];
    assign NewCRC[2] = D[46] ^ D[44] ^ D[43] ^ D[42] ^ D[41] ^ D[39] ^ D[38] ^ 
                D[34] ^ D[32] ^ D[30] ^ D[28] ^ D[27] ^ D[24] ^ D[22] ^ 
                D[19] ^ D[14] ^ D[13] ^ D[10] ^ D[9] ^ D[7] ^ D[6] ^ 
                D[5] ^ D[2] ^ D[1] ^ D[0];
    assign NewCRC[3] = D[47] ^ D[45] ^ D[44] ^ D[43] ^ D[42] ^ D[40] ^ D[39] ^ 
                D[35] ^ D[33] ^ D[31] ^ D[29] ^ D[28] ^ D[25] ^ D[23] ^ 
                D[20] ^ D[15] ^ D[14] ^ D[11] ^ D[10] ^ D[8] ^ D[7] ^ 
                D[6] ^ D[3] ^ D[2] ^ D[1];
    assign NewCRC[4] = D[45] ^ D[44] ^ D[43] ^ D[42] ^ D[40] ^ D[37] ^ D[35] ^ 
                D[33] ^ D[32] ^ D[31] ^ D[27] ^ D[21] ^ D[20] ^ D[18] ^ 
                D[17] ^ D[14] ^ D[13] ^ D[12] ^ D[11] ^ D[9] ^ D[6] ^ 
                D[4] ^ D[2] ^ D[1] ^ D[0];
    assign NewCRC[5] = D[46] ^ D[45] ^ D[44] ^ D[43] ^ D[41] ^ D[38] ^ D[36] ^ 
                D[34] ^ D[33] ^ D[32] ^ D[28] ^ D[22] ^ D[21] ^ D[19] ^ 
                D[18] ^ D[15] ^ D[14] ^ D[13] ^ D[12] ^ D[10] ^ D[7] ^ 
                D[5] ^ D[3] ^ D[2] ^ D[1];
    assign NewCRC[6] = D[47] ^ D[45] ^ D[44] ^ D[41] ^ D[39] ^ D[36] ^ D[31] ^ 
                D[30] ^ D[27] ^ D[26] ^ D[24] ^ D[23] ^ D[22] ^ D[19] ^ 
                D[18] ^ D[17] ^ D[11] ^ D[7] ^ D[4] ^ D[2] ^ D[1] ^ 
                D[0];
    assign NewCRC[7] = D[45] ^ D[41] ^ D[40] ^ D[36] ^ D[35] ^ D[34] ^ D[33] ^ 
                D[32] ^ D[30] ^ D[29] ^ D[28] ^ D[26] ^ D[25] ^ D[23] ^ 
                D[19] ^ D[17] ^ D[16] ^ D[15] ^ D[14] ^ D[13] ^ D[12] ^ 
                D[7] ^ D[6] ^ D[5] ^ D[2] ^ D[0];
					 
endmodule
