

module xor_32(
	input [31:0] a, input [31:0] b,
	output [31:0] out );

	assign out[0] 	=  a[0]  ^  b[0]; 
	assign out[1] 	=  a[1]  ^  b[1]; 
	assign out[2] 	=  a[2]  ^  b[2]; 
	assign out[3] 	=  a[3]  ^  b[3]; 
	assign out[4] 	=  a[4]  ^  b[4]; 
	assign out[5] 	=  a[5]  ^  b[5]; 
	assign out[6] 	=  a[6]  ^  b[6]; 
	assign out[7] 	=  a[7]  ^  b[7]; 
	assign out[8] 	=  a[8]  ^  b[8]; 
	assign out[9] 	=  a[9]  ^  b[9]; 
	assign out[10]	=  a[10] ^  b[10]; 
	assign out[11] 	=  a[11] ^  b[11]; 
	assign out[12] 	=  a[12] ^  b[12]; 
	assign out[13] 	=  a[13] ^  b[13]; 
	assign out[14] 	=  a[14] ^  b[14]; 
	assign out[15] 	=  a[15] ^  b[15]; 
	assign out[16] 	=  a[16] ^  b[16]; 
	assign out[17] 	=  a[17] ^  b[17]; 
	assign out[18] 	=  a[18] ^  b[18]; 
	assign out[19] 	=  a[19] ^  b[19]; 
	assign out[20] 	=  a[20] ^  b[20]; 
	assign out[21] 	=  a[21] ^  b[21]; 
	assign out[22] 	=  a[22] ^  b[22]; 
	assign out[23] 	=  a[23] ^  b[23];
	assign out[24] 	=  a[24] ^  b[24]; 
	assign out[25]	=  a[25] ^  b[25]; 
	assign out[26] 	=  a[26] ^  b[26]; 
	assign out[27] 	=  a[27] ^  b[27]; 
	assign out[28] 	=  a[28] ^  b[28]; 
	assign out[29] 	=  a[29] ^  b[29]; 
	assign out[30] 	=  a[30] ^  b[30];
	assign out[31] 	=  a[31] ^  b[31];
endmodule
