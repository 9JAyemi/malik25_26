
module full_adder (
    input a,
    input b,
    input cin,
    output sum,
    output cout
);

    assign sum = a ^ b ^ cin;
    assign cout = (a & b) | (a & cin) | (b & cin);

endmodule

module four_bit_adder (
    input [3:0] a,
    input [3:0] b,
    output [3:0] sum,
    output cout
);

    wire [2:0] c;

    full_adder fa1(a[0], b[0], 1'b0, sum[0], c[0]);
    full_adder fa2(a[1], b[1], c[0], sum[1], c[1]);
    full_adder fa3(a[2], b[2], c[1], sum[2], c[2]);
    full_adder fa4(a[3], b[3], c[2], sum[3], cout);

endmodule

module top_module (
    input [3:0] a,
    input [3:0] b,
    output [4:0] sum
);

    wire [2:0] c;

    four_bit_adder fa(a, b, sum[3:0], c[2]);
    assign sum[4] = c[2];

endmodule
