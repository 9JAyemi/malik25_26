
module muxed_ctrl_data(
  input [5:0] ByteCnt,
  input DlyCrcEn,
  input [1:0] DlyCrcCnt,
  input [47:0] MAC,
  input [15:0] TxPauseTV,
  input MTxClk,
  input TxReset,
  output reg [7:0] ControlData
);

reg [7:0] MuxedCtrlData;

always @ (ByteCnt or DlyCrcEn or MAC or TxPauseTV or DlyCrcCnt) begin
  case(ByteCnt)
    6'h0: if(~DlyCrcEn | DlyCrcEn & (&DlyCrcCnt[1:0]))
           MuxedCtrlData[7:0] = 8'h01; // Reserved Multicast Address
         else
           MuxedCtrlData[7:0] = 8'h0;
    6'h2: MuxedCtrlData[7:0] = 8'h80;
    6'h4: MuxedCtrlData[7:0] = 8'hC2;
    6'h6: MuxedCtrlData[7:0] = 8'h00;
    6'h8: MuxedCtrlData[7:0] = 8'h00;
    6'hA: MuxedCtrlData[7:0] = 8'h01;
    6'hC: MuxedCtrlData[7:0] = MAC[47:40];
    6'hE: MuxedCtrlData[7:0] = MAC[39:32];
    6'h10: MuxedCtrlData[7:0] = MAC[31:24];
    6'h12: MuxedCtrlData[7:0] = MAC[23:16];
    6'h14: MuxedCtrlData[7:0] = MAC[15:8];
    6'h16: MuxedCtrlData[7:0] = MAC[7:0];
    6'h18: MuxedCtrlData[7:0] = 8'h88; // Type/Length
    6'h1A: MuxedCtrlData[7:0] = 8'h08;
    6'h1C: MuxedCtrlData[7:0] = 8'h00; // Opcode
    6'h1E: MuxedCtrlData[7:0] = 8'h01;
    6'h20: MuxedCtrlData[7:0] = TxPauseTV[15:8]; // Pause timer value
    6'h22: MuxedCtrlData[7:0] = TxPauseTV[7:0];
    default: MuxedCtrlData[7:0] = 8'h0;
  endcase
end

always @ (posedge MTxClk or posedge TxReset) begin
  if(TxReset)
    ControlData[7:0] <= 8'h0;
  else if(~ByteCnt[0])
    ControlData[7:0] <= MuxedCtrlData[7:0];
end

endmodule