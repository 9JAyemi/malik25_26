
module my_inverter (
    output Y, // output
    input  A  // input
);

    not (Y, A);
endmodule