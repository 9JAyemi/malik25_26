module ay_note_ram(addr, data);
input wire [6:0] addr;
output wire [11:0] data; reg [11:0] note_ram [0:127];
initial begin
  note_ram[0] <= 12'd03977;
  note_ram[1] <= 12'd03977;
  note_ram[2] <= 12'd03977;
  note_ram[3] <= 12'd03977;
  note_ram[4] <= 12'd03977;
  note_ram[5] <= 12'd03977;
  note_ram[6] <= 12'd03977;
  note_ram[7] <= 12'd03977;
  note_ram[8] <= 12'd03977;
  note_ram[9] <= 12'd03977;
  note_ram[10] <= 12'd03977;
  note_ram[11] <= 12'd03977;
  note_ram[12] <= 12'd03977;
  note_ram[13] <= 12'd03977;
  note_ram[14] <= 12'd03977;
  note_ram[15] <= 12'd03977;
  note_ram[16] <= 12'd03977;
  note_ram[17] <= 12'd03977;
  note_ram[18] <= 12'd03977;
  note_ram[19] <= 12'd03977;
  note_ram[20] <= 12'd03977;
  note_ram[21] <= 12'd03977;
  note_ram[22] <= 12'd03754;
  note_ram[23] <= 12'd03543;
  note_ram[24] <= 12'd03344;
  note_ram[25] <= 12'd03157;
  note_ram[26] <= 12'd02980;
  note_ram[27] <= 12'd02812;
  note_ram[28] <= 12'd02655;
  note_ram[29] <= 12'd02506;
  note_ram[30] <= 12'd02365;
  note_ram[31] <= 12'd02232;
  note_ram[32] <= 12'd02107;
  note_ram[33] <= 12'd01989;
  note_ram[34] <= 12'd01877;
  note_ram[35] <= 12'd01772;
  note_ram[36] <= 12'd01672;
  note_ram[37] <= 12'd01578;
  note_ram[38] <= 12'd01490;
  note_ram[39] <= 12'd01406;
  note_ram[40] <= 12'd01327;
  note_ram[41] <= 12'd01253;
  note_ram[42] <= 12'd01182;
  note_ram[43] <= 12'd01116;
  note_ram[44] <= 12'd01053;
  note_ram[45] <= 12'd0994;
  note_ram[46] <= 12'd0939;
  note_ram[47] <= 12'd0886;
  note_ram[48] <= 12'd0836;
  note_ram[49] <= 12'd0789;
  note_ram[50] <= 12'd0745;
  note_ram[51] <= 12'd0703;
  note_ram[52] <= 12'd0664;
  note_ram[53] <= 12'd0626;
  note_ram[54] <= 12'd0591;
  note_ram[55] <= 12'd0558;
  note_ram[56] <= 12'd0527;
  note_ram[57] <= 12'd0497;
  note_ram[58] <= 12'd0469;
  note_ram[59] <= 12'd0443;
  note_ram[60] <= 12'd0418;
  note_ram[61] <= 12'd0395;
  note_ram[62] <= 12'd0372;
  note_ram[63] <= 12'd0352;
  note_ram[64] <= 12'd0332;
  note_ram[65] <= 12'd0313;
  note_ram[66] <= 12'd0296;
  note_ram[67] <= 12'd0279;
  note_ram[68] <= 12'd0263;
  note_ram[69] <= 12'd0249;
  note_ram[70] <= 12'd0235;
  note_ram[71] <= 12'd0221;
  note_ram[72] <= 12'd0209;
  note_ram[73] <= 12'd0197;
  note_ram[74] <= 12'd0186;
  note_ram[75] <= 12'd0176;
  note_ram[76] <= 12'd0166;
  note_ram[77] <= 12'd0157;
  note_ram[78] <= 12'd0148;
  note_ram[79] <= 12'd0140;
  note_ram[80] <= 12'd0132;
  note_ram[81] <= 12'd0124;
  note_ram[82] <= 12'd0117;
  note_ram[83] <= 12'd0111;
  note_ram[84] <= 12'd0105;
  note_ram[85] <= 12'd099;
  note_ram[86] <= 12'd093;
  note_ram[87] <= 12'd088;
  note_ram[88] <= 12'd083;
  note_ram[89] <= 12'd078;
  note_ram[90] <= 12'd074;
  note_ram[91] <= 12'd070;
  note_ram[92] <= 12'd066;
  note_ram[93] <= 12'd062;
  note_ram[94] <= 12'd059;
  note_ram[95] <= 12'd055;
  note_ram[96] <= 12'd052;
  note_ram[97] <= 12'd049;
  note_ram[98] <= 12'd047;
  note_ram[99] <= 12'd044;
  note_ram[100] <= 12'd041;
  note_ram[101] <= 12'd039;
  note_ram[102] <= 12'd037;
  note_ram[103] <= 12'd035;
  note_ram[104] <= 12'd033;
  note_ram[105] <= 12'd031;
  note_ram[106] <= 12'd029;
  note_ram[107] <= 12'd028;
  note_ram[108] <= 12'd026;
  note_ram[109] <= 12'd025;
  note_ram[110] <= 12'd023;
  note_ram[111] <= 12'd022;
  note_ram[112] <= 12'd021;
  note_ram[113] <= 12'd020;
  note_ram[114] <= 12'd018;
  note_ram[115] <= 12'd017;
  note_ram[116] <= 12'd016;
  note_ram[117] <= 12'd016;
  note_ram[118] <= 12'd015;
  note_ram[119] <= 12'd014;
  note_ram[120] <= 12'd013;
  note_ram[121] <= 12'd012;
  note_ram[122] <= 12'd012;
  note_ram[123] <= 12'd011;
  note_ram[124] <= 12'd010;
  note_ram[125] <= 12'd010;
  note_ram[126] <= 12'd09;
  note_ram[127] <= 12'd09;
end

assign data = note_ram[addr];

endmodule
