// SVA checker for bpm_from_interval
// Binds a golden lookup and concise assertions + coverage.

module bpm_from_interval_sva (
  input logic [31:0] counter,
  input logic [7:0]  default_bpm,
  input logic [7:0]  counted_bpm
);

  function automatic byte unsigned ref_bpm(input logic [31:0] counter_i, input byte unsigned dflt);
    `define STEP(T,V) else if (counter_i < 32'd``T) return 8'd``V;
    if (counter_i < 32'd23529) return 8'd254;
    `STEP(23622,253)
    `STEP(23715,252)
    `STEP(23809,251)
    `STEP(23904,250)
    `STEP(24000,249)
    `STEP(24096,248)
    `STEP(24193,247)
    `STEP(24291,246)
    `STEP(24390,245)
    `STEP(24489,244)
    `STEP(24590,243)
    `STEP(24691,242)
    `STEP(24793,241)
    `STEP(24896,240)
    `STEP(25000,239)
    `STEP(25104,238)
    `STEP(25210,237)
    `STEP(25316,236)
    `STEP(25423,235)
    `STEP(25531,234)
    `STEP(25641,233)
    `STEP(25751,232)
    `STEP(25862,231)
    `STEP(25974,230)
    `STEP(26086,229)
    `STEP(26200,228)
    `STEP(26315,227)
    `STEP(26431,226)
    `STEP(26548,225)
    `STEP(26666,224)
    `STEP(26785,223)
    `STEP(26905,222)
    `STEP(27027,221)
    `STEP(27149,220)
    `STEP(27272,219)
    `STEP(27397,218)
    `STEP(27522,217)
    `STEP(27649,216)
    `STEP(27777,215)
    `STEP(27906,214)
    `STEP(28037,213)
    `STEP(28169,212)
    `STEP(28301,211)
    `STEP(28436,210)
    `STEP(28571,209)
    `STEP(28708,208)
    `STEP(28846,207)
    `STEP(28985,206)
    `STEP(29126,205)
    `STEP(29268,204)
    `STEP(29411,203)
    `STEP(29556,202)
    `STEP(29702,201)
    `STEP(29850,200)
    `STEP(30000,199)
    `STEP(30150,198)
    `STEP(30303,197)
    `STEP(30456,196)
    `STEP(30612,195)
    `STEP(30769,194)
    `STEP(30927,193)
    `STEP(31088,192)
    `STEP(31250,191)
    `STEP(31413,190)
    `STEP(31578,189)
    `STEP(31746,188)
    `STEP(31914,187)
    `STEP(32085,186)
    `STEP(32258,185)
    `STEP(32432,184)
    `STEP(32608,183)
    `STEP(32786,182)
    `STEP(32967,181)
    `STEP(33149,180)
    `STEP(33333,179)
    `STEP(33519,178)
    `STEP(33707,177)
    `STEP(33898,176)
    `STEP(34090,175)
    `STEP(34285,174)
    `STEP(34482,173)
    `STEP(34682,172)
    `STEP(34883,171)
    `STEP(35087,170)
    `STEP(35294,169)
    `STEP(35502,168)
    `STEP(35714,167)
    `STEP(35928,166)
    `STEP(36144,165)
    `STEP(36363,164)
    `STEP(36585,163)
    `STEP(36809,162)
    `STEP(37037,161)
    `STEP(37267,160)
    `STEP(37500,159)
    `STEP(37735,158)
    `STEP(37974,157)
    `STEP(38216,156)
    `STEP(38461,155)
    `STEP(38709,154)
    `STEP(38961,153)
    `STEP(39215,152)
    `STEP(39473,151)
    `STEP(39735,150)
    `STEP(40000,149)
    `STEP(40268,148)
    `STEP(40540,147)
    `STEP(40816,146)
    `STEP(41095,145)
    `STEP(41379,144)
    `STEP(41666,143)
    `STEP(41958,142)
    `STEP(42253,141)
    `STEP(42553,140)
    `STEP(42857,139)
    `STEP(43165,138)
    `STEP(43478,137)
    `STEP(43795,136)
    `STEP(44117,135)
    `STEP(44444,134)
    `STEP(44776,133)
    `STEP(45112,132)
    `STEP(45454,131)
    `STEP(45801,130)
    `STEP(46153,129)
    `STEP(46511,128)
    `STEP(46875,127)
    `STEP(47244,126)
    `STEP(47619,125)
    `STEP(48000,124)
    `STEP(48387,123)
    `STEP(48780,122)
    `STEP(49180,121)
    `STEP(49586,120)
    `STEP(50000,119)
    `STEP(50420,118)
    `STEP(50847,117)
    `STEP(51282,116)
    `STEP(51724,115)
    `STEP(52173,114)
    `STEP(52631,113)
    `STEP(53097,112)
    `STEP(53571,111)
    `STEP(54054,110)
    `STEP(54545,109)
    `STEP(55045,108)
    `STEP(55555,107)
    `STEP(56074,106)
    `STEP(56603,105)
    `STEP(57142,104)
    `STEP(57692,103)
    `STEP(58252,102)
    `STEP(58823,101)
    `STEP(59405,100)
    `STEP(60000,99)
    `STEP(60606,98)
    `STEP(61224,97)
    `STEP(61855,96)
    `STEP(62500,95)
    `STEP(63157,94)
    `STEP(63829,93)
    `STEP(64516,92)
    `STEP(65217,91)
    `STEP(65934,90)
    `STEP(66666,89)
    `STEP(67415,88)
    `STEP(68181,87)
    `STEP(68965,86)
    `STEP(69767,85)
    `STEP(70588,84)
    `STEP(71428,83)
    `STEP(72289,82)
    `STEP(73170,81)
    `STEP(74074,80)
    `STEP(75000,79)
    `STEP(75949,78)
    `STEP(76923,77)
    `STEP(77922,76)
    `STEP(78947,75)
    `STEP(80000,74)
    `STEP(81081,73)
    `STEP(82191,72)
    `STEP(83333,71)
    `STEP(84507,70)
    `STEP(85714,69)
    `STEP(86956,68)
    `STEP(88235,67)
    `STEP(89552,66)
    `STEP(90909,65)
    `STEP(92307,64)
    `STEP(93750,63)
    `STEP(95238,62)
    `STEP(96774,61)
    `STEP(98360,60)
    `STEP(100000,59)
    `STEP(101694,58)
    `STEP(103448,57)
    `STEP(105263,56)
    `STEP(107142,55)
    `STEP(109090,54)
    `STEP(111111,53)
    `STEP(113207,52)
    `STEP(115384,51)
    `STEP(117647,50)
    `STEP(120000,49)
    `STEP(122448,48)
    `STEP(125000,47)
    `STEP(127659,46)
    `STEP(130434,45)
    `STEP(133333,44)
    `STEP(136363,43)
    `STEP(139534,42)
    `STEP(142857,41)
    `STEP(146341,40)
    `STEP(150000,39)
    `STEP(153846,38)
    `STEP(157894,37)
    `STEP(162162,36)
    `STEP(166666,35)
    `STEP(171428,34)
    `STEP(176470,33)
    `STEP(181818,32)
    `STEP(187500,31)
    `STEP(193548,30)
    else return dflt;
    `undef STEP
  endfunction

  // Functional equivalence (combinational immediate SVA)
  always_comb begin
    byte unsigned exp = ref_bpm(counter, default_bpm);
    assert (counted_bpm === exp)
      else $error("bpm_from_interval: mismatch exp=%0d got=%0d counter=%0d default=%0d",
                  exp, counted_bpm, counter, default_bpm);

    if (!$isunknown({counter, default_bpm}))
      assert (!$isunknown(counted_bpm))
        else $error("bpm_from_interval: X/Z on counted_bpm");

    if (counted_bpm !== default_bpm)
      assert (counted_bpm inside {[8'd30:8'd254]})
        else $error("bpm_from_interval: out-of-range LUT value %0d", counted_bpm);

    if (counter >= 32'd193548)
      assert (counted_bpm == default_bpm)
        else $error("bpm_from_interval: default path violated");
  end

  // Coverage
  covergroup cg_bpm @(counter or default_bpm or counted_bpm);
    cp_val: coverpoint counted_bpm {
      bins lut_vals[] = {[8'd30:8'd254]};
    }
    cp_default_used: coverpoint (counted_bpm == default_bpm) iff (counter >= 32'd193548) {
      bins used = {1};
    }
    cp_edges: coverpoint counter {
      bins first_minus = {32'd23528};
      bins first_edge  = {32'd23529};
      bins last_minus  = {32'd193547};
      bins last_edge   = {32'd193548};
    }
  endgroup
  cg_bpm cg = new();

endmodule

bind bpm_from_interval bpm_from_interval_sva bpm_from_interval_sva_i (
  .counter(counter),
  .default_bpm(default_bpm),
  .counted_bpm(counted_bpm)
);