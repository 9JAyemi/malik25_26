
module nor4_gate(
    input A,
    input B,
    input C,
    input D,
    output Y
);

    nor (Y, A, B, C, D);

endmodule
