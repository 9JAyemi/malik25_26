

module bpm_from_interval(
    input [31:0] counter, 			  input wire [7:0] default_bpm,  output wire [7:0] counted_bpm  );
								
	assign counted_bpm = (counter < 32'd23529 ) ? 254 : (counter < 32'd23622 ) ? 253 : (counter < 32'd23715 ) ? 252 : (counter < 32'd23809 ) ? 251 : 
								(counter < 32'd23904 ) ? 250 :
								(counter < 32'd24000 ) ? 249 :
								(counter < 32'd24096 ) ? 248 :
								(counter < 32'd24193 ) ? 247 :
								(counter < 32'd24291 ) ? 246 :
								(counter < 32'd24390 ) ? 245 :
								(counter < 32'd24489 ) ? 244 :
								(counter < 32'd24590 ) ? 243 :
								(counter < 32'd24691 ) ? 242 :
								(counter < 32'd24793 ) ? 241 :
								(counter < 32'd24896 ) ? 240 :
								(counter < 32'd25000 ) ? 239 :
								(counter < 32'd25104 ) ? 238 :
								(counter < 32'd25210 ) ? 237 :
								(counter < 32'd25316 ) ? 236 :
								(counter < 32'd25423 ) ? 235 :
								(counter < 32'd25531 ) ? 234 :
								(counter < 32'd25641 ) ? 233 :
								(counter < 32'd25751 ) ? 232 :
								(counter < 32'd25862 ) ? 231 :
								(counter < 32'd25974 ) ? 230 :
								(counter < 32'd26086 ) ? 229 :
								(counter < 32'd26200 ) ? 228 :
								(counter < 32'd26315 ) ? 227 :
								(counter < 32'd26431 ) ? 226 :
								(counter < 32'd26548 ) ? 225 :
								(counter < 32'd26666 ) ? 224 :
								(counter < 32'd26785 ) ? 223 :
								(counter < 32'd26905 ) ? 222 :
								(counter < 32'd27027 ) ? 221 :
								(counter < 32'd27149 ) ? 220 :
								(counter < 32'd27272 ) ? 219 :
								(counter < 32'd27397 ) ? 218 :
								(counter < 32'd27522 ) ? 217 :
								(counter < 32'd27649 ) ? 216 :
								(counter < 32'd27777 ) ? 215 :
								(counter < 32'd27906 ) ? 214 :
								(counter < 32'd28037 ) ? 213 :
								(counter < 32'd28169 ) ? 212 :
								(counter < 32'd28301 ) ? 211 :
								(counter < 32'd28436 ) ? 210 :
								(counter < 32'd28571 ) ? 209 :
								(counter < 32'd28708 ) ? 208 :
								(counter < 32'd28846 ) ? 207 :
								(counter < 32'd28985 ) ? 206 :
								(counter < 32'd29126 ) ? 205 :
								(counter < 32'd29268 ) ? 204 :
								(counter < 32'd29411 ) ? 203 :
								(counter < 32'd29556 ) ? 202 :
								(counter < 32'd29702 ) ? 201 :
								(counter < 32'd29850 ) ? 200 :
								(counter < 32'd30000 ) ? 199 :
								(counter < 32'd30150 ) ? 198 :
								(counter < 32'd30303 ) ? 197 :
								(counter < 32'd30456 ) ? 196 :
								(counter < 32'd30612 ) ? 195 :
								(counter < 32'd30769 ) ? 194 :
								(counter < 32'd30927 ) ? 193 :
								(counter < 32'd31088 ) ? 192 :
								(counter < 32'd31250 ) ? 191 :
								(counter < 32'd31413 ) ? 190 :
								(counter < 32'd31578 ) ? 189 :
								(counter < 32'd31746 ) ? 188 :
								(counter < 32'd31914 ) ? 187 :
								(counter < 32'd32085 ) ? 186 :
								(counter < 32'd32258 ) ? 185 :
								(counter < 32'd32432 ) ? 184 :
								(counter < 32'd32608 ) ? 183 :
								(counter < 32'd32786 ) ? 182 :
								(counter < 32'd32967 ) ? 181 :
								(counter < 32'd33149 ) ? 180 :
								(counter < 32'd33333 ) ? 179 :
								(counter < 32'd33519 ) ? 178 :
								(counter < 32'd33707 ) ? 177 :
								(counter < 32'd33898 ) ? 176 :
								(counter < 32'd34090 ) ? 175 :
								(counter < 32'd34285 ) ? 174 :
								(counter < 32'd34482 ) ? 173 :
								(counter < 32'd34682 ) ? 172 :
								(counter < 32'd34883 ) ? 171 :
								(counter < 32'd35087 ) ? 170 :
								(counter < 32'd35294 ) ? 169 :
								(counter < 32'd35502 ) ? 168 :
								(counter < 32'd35714 ) ? 167 :
								(counter < 32'd35928 ) ? 166 :
								(counter < 32'd36144 ) ? 165 :
								(counter < 32'd36363 ) ? 164 :
								(counter < 32'd36585 ) ? 163 :
								(counter < 32'd36809 ) ? 162 :
								(counter < 32'd37037 ) ? 161 :
								(counter < 32'd37267 ) ? 160 :
								(counter < 32'd37500 ) ? 159 :
								(counter < 32'd37735 ) ? 158 :
								(counter < 32'd37974 ) ? 157 :
								(counter < 32'd38216 ) ? 156 :
								(counter < 32'd38461 ) ? 155 :
								(counter < 32'd38709 ) ? 154 :
								(counter < 32'd38961 ) ? 153 :
								(counter < 32'd39215 ) ? 152 :
								(counter < 32'd39473 ) ? 151 :
								(counter < 32'd39735 ) ? 150 :
								(counter < 32'd40000 ) ? 149 :
								(counter < 32'd40268 ) ? 148 :
								(counter < 32'd40540 ) ? 147 :
								(counter < 32'd40816 ) ? 146 :
								(counter < 32'd41095 ) ? 145 :
								(counter < 32'd41379 ) ? 144 :
								(counter < 32'd41666 ) ? 143 :
								(counter < 32'd41958 ) ? 142 :
								(counter < 32'd42253 ) ? 141 :
								(counter < 32'd42553 ) ? 140 :
								(counter < 32'd42857 ) ? 139 :
								(counter < 32'd43165 ) ? 138 :
								(counter < 32'd43478 ) ? 137 :
								(counter < 32'd43795 ) ? 136 :
								(counter < 32'd44117 ) ? 135 :
								(counter < 32'd44444 ) ? 134 :
								(counter < 32'd44776 ) ? 133 :
								(counter < 32'd45112 ) ? 132 :
								(counter < 32'd45454 ) ? 131 :
								(counter < 32'd45801 ) ? 130 :
								(counter < 32'd46153 ) ? 129 :
								(counter < 32'd46511 ) ? 128 :
								(counter < 32'd46875 ) ? 127 :
								(counter < 32'd47244 ) ? 126 :
								(counter < 32'd47619 ) ? 125 :
								(counter < 32'd48000 ) ? 124 :
								(counter < 32'd48387 ) ? 123 :
								(counter < 32'd48780 ) ? 122 :
								(counter < 32'd49180 ) ? 121 :
								(counter < 32'd49586 ) ? 120 :
								(counter < 32'd50000 ) ? 119 :
								(counter < 32'd50420 ) ? 118 :
								(counter < 32'd50847 ) ? 117 :
								(counter < 32'd51282 ) ? 116 :
								(counter < 32'd51724 ) ? 115 :
								(counter < 32'd52173 ) ? 114 :
								(counter < 32'd52631 ) ? 113 :
								(counter < 32'd53097 ) ? 112 :
								(counter < 32'd53571 ) ? 111 :
								(counter < 32'd54054 ) ? 110 :
								(counter < 32'd54545 ) ? 109 :
								(counter < 32'd55045 ) ? 108 :
								(counter < 32'd55555 ) ? 107 :
								(counter < 32'd56074 ) ? 106 :
								(counter < 32'd56603 ) ? 105 :
								(counter < 32'd57142 ) ? 104 :
								(counter < 32'd57692 ) ? 103 :
								(counter < 32'd58252 ) ? 102 :
								(counter < 32'd58823 ) ? 101 :
								(counter < 32'd59405 ) ? 100 :
								(counter < 32'd60000 ) ? 99 :
								(counter < 32'd60606 ) ? 98 :
								(counter < 32'd61224 ) ? 97 :
								(counter < 32'd61855 ) ? 96 :
								(counter < 32'd62500 ) ? 95 :
								(counter < 32'd63157 ) ? 94 :
								(counter < 32'd63829 ) ? 93 :
								(counter < 32'd64516 ) ? 92 :
								(counter < 32'd65217 ) ? 91 :
								(counter < 32'd65934 ) ? 90 :
								(counter < 32'd66666 ) ? 89 :
								(counter < 32'd67415 ) ? 88 :
								(counter < 32'd68181 ) ? 87 :
								(counter < 32'd68965 ) ? 86 :
								(counter < 32'd69767 ) ? 85 :
								(counter < 32'd70588 ) ? 84 :
								(counter < 32'd71428 ) ? 83 :
								(counter < 32'd72289 ) ? 82 :
								(counter < 32'd73170 ) ? 81 :
								(counter < 32'd74074 ) ? 80 :
								(counter < 32'd75000 ) ? 79 :
								(counter < 32'd75949 ) ? 78 :
								(counter < 32'd76923 ) ? 77 :
								(counter < 32'd77922 ) ? 76 :
								(counter < 32'd78947 ) ? 75 :
								(counter < 32'd80000 ) ? 74 :
								(counter < 32'd81081 ) ? 73 :
								(counter < 32'd82191 ) ? 72 :
								(counter < 32'd83333 ) ? 71 :
								(counter < 32'd84507 ) ? 70 :
								(counter < 32'd85714 ) ? 69 :
								(counter < 32'd86956 ) ? 68 :
								(counter < 32'd88235 ) ? 67 :
								(counter < 32'd89552 ) ? 66 :
								(counter < 32'd90909 ) ? 65 :
								(counter < 32'd92307 ) ? 64 :
								(counter < 32'd93750 ) ? 63 :
								(counter < 32'd95238 ) ? 62 :
								(counter < 32'd96774 ) ? 61 :
								(counter < 32'd98360 ) ? 60 :
								(counter < 32'd100000 ) ? 59 :
								(counter < 32'd101694 ) ? 58 :
								(counter < 32'd103448 ) ? 57 :
								(counter < 32'd105263 ) ? 56 :
								(counter < 32'd107142 ) ? 55 :
								(counter < 32'd109090 ) ? 54 :
								(counter < 32'd111111 ) ? 53 :
								(counter < 32'd113207 ) ? 52 :
								(counter < 32'd115384 ) ? 51 :
								(counter < 32'd117647 ) ? 50 :
								(counter < 32'd120000 ) ? 49 :
								(counter < 32'd122448 ) ? 48 :
								(counter < 32'd125000 ) ? 47 :
								(counter < 32'd127659 ) ? 46 :
								(counter < 32'd130434 ) ? 45 :
								(counter < 32'd133333 ) ? 44 :
								(counter < 32'd136363 ) ? 43 :
								(counter < 32'd139534 ) ? 42 :
								(counter < 32'd142857 ) ? 41 :
								(counter < 32'd146341 ) ? 40 :
								(counter < 32'd150000 ) ? 39 :
								(counter < 32'd153846 ) ? 38 :
								(counter < 32'd157894 ) ? 37 :
								(counter < 32'd162162 ) ? 36 :
								(counter < 32'd166666 ) ? 35 :
								(counter < 32'd171428 ) ? 34 :
								(counter < 32'd176470 ) ? 33 :
								(counter < 32'd181818 ) ? 32 :
								(counter < 32'd187500 ) ? 31 :
								(counter < 32'd193548 ) ? 30 : default_bpm;
endmodule
