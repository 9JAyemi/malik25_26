
module sky130_fd_sc_hs__o21a_1 (A1, A2, B1, VPWR, VGND, Y);
  input A1, A2, B1, VPWR, VGND;
  output Y;

  // Implementation of the module

endmodule

module sky130_fd_sc_hs__o21a_2 (A1, A2, B1, VPWR, VGND, Y);
  input A1, A2, B1, VPWR, VGND;
  output Y;

  assign Y = (A1 & A2) | B1;

endmodule
