
module pll_lock_lookup(
    input clk,
    input [6:0] divider,
    output reg [39:0] value
    );
     reg [39:0] lookup [0:64];
    wire [5:0] addr;
   initial
   begin
            lookup[00]=40'b00110_00110_1111101000_1111101001_0000000001;
            lookup[01]=40'b00110_00110_1111101000_1111101001_0000000001;
            lookup[02]=40'b01000_01000_1111101000_1111101001_0000000001;
            lookup[03]=40'b01011_01011_1111101000_1111101001_0000000001;
            lookup[04]=40'b01110_01110_1111101000_1111101001_0000000001;
            lookup[05]=40'b10001_10001_1111101000_1111101001_0000000001;
            lookup[06]=40'b10011_10011_1111101000_1111101001_0000000001;
            lookup[07]=40'b10110_10110_1111101000_1111101001_0000000001;
            lookup[08]=40'b11001_11001_1111101000_1111101001_0000000001;
            lookup[09]=40'b11100_11100_1111101000_1111101001_0000000001;
            lookup[10]=40'b11111_11111_1110000100_1111101001_0000000001;
            lookup[11]=40'b11111_11111_1100111001_1111101001_0000000001;
            lookup[12]=40'b11111_11111_1011101110_1111101001_0000000001;
            lookup[13]=40'b11111_11111_1010111100_1111101001_0000000001;
            lookup[14]=40'b11111_11111_1010001010_1111101001_0000000001;
            lookup[15]=40'b11111_11111_1001110001_1111101001_0000000001;
            lookup[16]=40'b11111_11111_1000111111_1111101001_0000000001;
            lookup[17]=40'b11111_11111_1000100110_1111101001_0000000001;
            lookup[18]=40'b11111_11111_1000001101_1111101001_0000000001;
            lookup[19]=40'b11111_11111_0111110100_1111101001_0000000001;
            lookup[20]=40'b11111_11111_0111011011_1111101001_0000000001;
            lookup[21]=40'b11111_11111_0111000010_1111101001_0000000001;
            lookup[22]=40'b11111_11111_0110101001_1111101001_0000000001;
            lookup[23]=40'b11111_11111_0110010000_1111101001_0000000001;
            lookup[24]=40'b11111_11111_0110010000_1111101001_0000000001;
            lookup[25]=40'b11111_11111_0101110111_1111101001_0000000001;
            lookup[26]=40'b11111_11111_0101011110_1111101001_0000000001;
            lookup[27]=40'b11111_11111_0101011110_1111101001_0000000001;
            lookup[28]=40'b11111_11111_0101000101_1111101001_0000000001;
            lookup[29]=40'b11111_11111_0101000101_1111101001_0000000001;
            lookup[30]=40'b11111_11111_0100101100_1111101001_0000000001;
            lookup[31]=40'b11111_11111_0100101100_1111101001_0000000001;
            lookup[32]=40'b11111_11111_0100101100_1111101001_0000000001;
            lookup[33]=40'b11111_11111_0100010011_1111101001_0000000001;
            lookup[34]=40'b11111_11111_0100010011_1111101001_0000000001;
            lookup[35]=40'b11111_11111_0100010011_1111101001_0000000001;
            lookup[36]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[37]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[38]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[39]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[40]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[41]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[42]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[43]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[44]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[45]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[46]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[47]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[48]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[49]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[50]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[51]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[52]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[53]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[54]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[55]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[56]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[57]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[58]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[59]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[60]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[6]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[00]=40'b11111_11111_0011111010_1111101001_0000000001;
            lookup[00]=40'b11111_11111_0011111010_1111101001_0000000001;
   end
   
   assign addr = divider - 1;
   always @(posedge clk)
   begin
       value = lookup[addr];
   end 

endmodule
