module four_bit_adder(a, b, sum);
input [3:0] a;
input [3:0] b;
output [3:0] sum;

assign sum = a + b;

endmodule