module Vector(a, b, c);

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// I/O declarations

	
	input wire[1:0] a;

	
	input wire[1:0] b;

	
	output wire[1:0] c;

	////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	// The actual logic

	assign c = a & b;

endmodule