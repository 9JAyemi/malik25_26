module blinki (
  
  input Reset_n_i,
  
  input Clk_i,
  
  output reg LED_o,
  
  input[15:0] PeriodH_i,
  
  input[15:0] PeriodL_i
);

  localparam stStart   = 3'b000;
  localparam stOn      = 3'b001;
  localparam stOff     = 3'b010;
  reg  [2:0]             State;
  reg  [2:0]             NextState;
  reg                    TimerPreset;
  reg                    TimerEnable;
  wire                   TimerOvfl;

  always @(negedge Reset_n_i or posedge Clk_i)
  begin
    if (!Reset_n_i)
    begin
      State <= stStart;
    end
    else
    begin State <= NextState;
    end  
  end

  always @(State, TimerOvfl)
  begin  NextState     = State;
    TimerEnable   = 1'b1;
    TimerPreset   = 1'b0;
    case (State)
      stStart: begin
        TimerPreset   = 1'b1;
        NextState     = stOn;
      end
      stOn: begin
        LED_o = 1'b1;
        if (TimerOvfl == 1'b1)
        begin
          NextState     = stOff;
          TimerPreset   = 1'b1;
        end
      end
      stOff: begin
        LED_o = 1'b0;
        if (TimerOvfl == 1'b1)
        begin
          NextState     = stOn;
          TimerPreset   = 1'b1;
        end
      end
      default: begin
      end
    endcase
  end 

  reg [31:0] Timer;
  
  always @(negedge Reset_n_i or posedge Clk_i)
  begin
    if (!Reset_n_i)
    begin
      Timer <= 32'd0;
    end
    else
    begin
      if (TimerPreset)
      begin
        Timer <= {PeriodH_i, PeriodL_i};
      end
      else if (TimerEnable)
      begin
        Timer <= Timer - 1'b1;
      end
    end  
  end

  assign TimerOvfl = (Timer == 0) ? 1'b1 : 1'b0;

endmodule
