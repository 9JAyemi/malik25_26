module frame_rate (
    input inclk0,
    output reg c0,
    output reg c1,
    output reg locked
);

reg inclk0_d; // delayed inclk0 signal
reg locked_d; // delayed locked signal
reg locked_dd; // doubly delayed locked signal
reg c0_d; // delayed c0 signal
reg c1_d; // delayed c1 signal
reg c0_dd; // doubly delayed c0 signal
reg c1_dd; // doubly delayed c1 signal
reg locked_next; // next value of locked signal
reg c0_next; // next value of c0 signal
reg c1_next; // next value of c1 signal

parameter COUNT_MAX = 2; // number of clock cycles to wait before updating output signals

integer count = 0; // counter for number of clock cycles elapsed

always @(posedge inclk0)
begin
    // update delayed signals
    inclk0_d <= inclk0;
    c0_d <= c0_next;
    c1_d <= c1_next;
    locked_d <= locked_next;

    // update doubly delayed signals
    c0_dd <= c0_d;
    c1_dd <= c1_d;
    locked_dd <= locked_d;

    // update output signals
    if (count == COUNT_MAX)
    begin
        c0 <= c0_d;
        c1 <= c1_d;
        locked <= locked_d;

        // calculate next values of output signals
        c0_next <= ~c0_dd;
        c1_next <= c0_dd;
        locked_next <= (inclk0_d == locked_dd) ? 1 : 0;

        count <= 0;
    end
    else
    begin
        count <= count + 1;
    end
end

endmodule