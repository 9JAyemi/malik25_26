module top_module(
    input [2:0] sel,
    input [3:0] data0,
    input [3:0] data1,
    input [3:0] data2,
    input [3:0] data3,
    input [3:0] data4,
    input [3:0] data5,
    input [3:0] data6,
    input [3:0] data7,
    output [3:0] out
);

// 8-to-1 MUX implementation
assign out = (sel == 3'd0) ? data0 :
             (sel == 3'd1) ? data1 :
             (sel == 3'd2) ? data2 :
             (sel == 3'd3) ? data3 :
             (sel == 3'd4) ? data4 :
             (sel == 3'd5) ? data5 :
             (sel == 3'd6) ? data6 :
                             data7;

endmodule