
module channel_bridge (
    input clk,
    input reset_n,
    input in_valid,
    input [7:0] in_data,
    input [7:0] in_channel,
    input in_startofpacket,
    input in_endofpacket,
    output reg out_valid,
    output reg [7:0] out_data,
    output reg [7:0] out_channel,
    output reg out_startofpacket,
    output reg out_endofpacket
);

    reg [7:0] stored_data;
    reg [7:0] stored_channel;
    reg stored_startofpacket;
    reg stored_endofpacket;

    always @(posedge clk) begin
        if (!reset_n) begin
            out_valid <= 1'b0;
            out_data <= 8'd0;
            out_channel <= 8'd0;
            out_startofpacket <= 1'b0;
            out_endofpacket <= 1'b0;
        end else begin
            if (in_valid) begin
                stored_data <= in_data;
                stored_channel <= in_channel;
                stored_startofpacket <= in_startofpacket;
                stored_endofpacket <= in_endofpacket;
            end

            if (out_valid) begin
                out_data <= stored_data;
                out_channel <= stored_channel;
                out_startofpacket <= stored_startofpacket;
                out_endofpacket <= stored_endofpacket;

                if (in_channel > 8'd0) begin
                    out_valid <= 1'b0;
                    //$display("Simulation Message: Channel %d is suppressed", in_channel);
                end
            end else begin
                out_valid <= 1'b1;
            end
        end
    end

endmodule