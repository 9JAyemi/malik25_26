module xor_gate (
    input A,
    input B,
    output X
);

    assign X = A ^ B;

endmodule