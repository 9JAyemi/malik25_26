module decoder_4to16 (
    input [3:0] ABCD,
    output reg [15:0] Y
);

always @(*) begin
    case (ABCD)
        4'b0000: Y = 16'b1111_1111_1111_1110;
        4'b0001: Y = 16'b1111_1111_1111_1101;
        4'b0010: Y = 16'b1111_1111_1111_1011;
        4'b0011: Y = 16'b1111_1111_1111_0111;
        4'b0100: Y = 16'b1111_1111_1110_1111;
        4'b0101: Y = 16'b1111_1111_1101_1111;
        4'b0110: Y = 16'b1111_1111_1011_1111;
        4'b0111: Y = 16'b1111_1111_0111_1111;
        4'b1000: Y = 16'b1111_1110_1111_1111;
        4'b1001: Y = 16'b1111_1101_1111_1111;
        4'b1010: Y = 16'b1111_1011_1111_1111;
        4'b1011: Y = 16'b1111_0111_1111_1111;
        4'b1100: Y = 16'b1110_1111_1111_1111;
        4'b1101: Y = 16'b1101_1111_1111_1111;
        4'b1110: Y = 16'b1011_1111_1111_1111;
        4'b1111: Y = 16'b0111_1111_1111_1111;
        default: Y = 16'b1111_1111_1111_1111;
    endcase
end

endmodule