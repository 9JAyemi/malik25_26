module decoder_4to16 (
    input A,
    input B,
    input C,
    input D,
    output reg [15:0] Y
);

always @(*) begin
    if (A == 0 && B == 0 && C == 0 && D == 0) Y = 16'b1111111111111110;
    else if (A == 0 && B == 0 && C == 0 && D == 1) Y = 16'b1111111111111101;
    else if (A == 0 && B == 0 && C == 1 && D == 0) Y = 16'b1111111111111011;
    else if (A == 0 && B == 0 && C == 1 && D == 1) Y = 16'b1111111111110111;
    else if (A == 0 && B == 1 && C == 0 && D == 0) Y = 16'b1111111111101111;
    else if (A == 0 && B == 1 && C == 0 && D == 1) Y = 16'b1111111111011111;
    else if (A == 0 && B == 1 && C == 1 && D == 0) Y = 16'b1111111110111111;
    else if (A == 0 && B == 1 && C == 1 && D == 1) Y = 16'b1111111101111111;
    else if (A == 1 && B == 0 && C == 0 && D == 0) Y = 16'b1111111011111111;
    else if (A == 1 && B == 0 && C == 0 && D == 1) Y = 16'b1111110111111111;
    else if (A == 1 && B == 0 && C == 1 && D == 0) Y = 16'b1111101111111111;
    else if (A == 1 && B == 0 && C == 1 && D == 1) Y = 16'b1111011111111111;
    else if (A == 1 && B == 1 && C == 0 && D == 0) Y = 16'b1110111111111111;
    else if (A == 1 && B == 1 && C == 0 && D == 1) Y = 16'b1101111111111111;
    else if (A == 1 && B == 1 && C == 1 && D == 0) Y = 16'b1011111111111111;
    else if (A == 1 && B == 1 && C == 1 && D == 1) Y = 16'b0111111111111111;
end

endmodule