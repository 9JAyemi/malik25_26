module vga(input vclock,
            output reg [9:0] hcount,  // pixel number on current line
            output reg [9:0] vcount,  // line number
            output reg vsync,hsync,blank);

// VGA (640x480) @ 60 Hz
parameter VGA_HBLANKON  =  10'd639;
parameter VGA_HSYNCON   =  10'd655;
parameter VGA_HSYNCOFF  =  10'd751;
parameter VGA_HRESET    =  10'd799;
parameter VGA_VBLANKON  =  10'd479;
parameter VGA_VSYNCON   =  10'd490;
parameter VGA_VSYNCOFF  =  10'd492;
parameter VGA_VRESET    =  10'd523;

reg hblank,vblank;
wire hsyncon,hsyncoff,hreset,hblankon;
assign hblankon = (hcount == VGA_HBLANKON);
assign hsyncon = (hcount == VGA_HSYNCON);
assign hsyncoff = (hcount == VGA_HSYNCOFF);
assign hreset = (hcount == VGA_HRESET);

wire vsyncon,vsyncoff,vreset,vblankon;
assign vblankon = hreset & (vcount == VGA_VBLANKON);
assign vsyncon = hreset & (vcount == VGA_VSYNCON);
assign vsyncoff = hreset & (vcount == VGA_VSYNCOFF);
assign vreset = hreset & (vcount == VGA_VRESET);

// sync and blanking
wire next_hblank,next_vblank;
assign next_hblank = hreset ? 0 : hblankon ? 1 : hblank;
assign next_vblank = vreset ? 0 : vblankon ? 1 : vblank;

// VGA controller
always @(posedge vclock) begin
    if (hcount == 799 && vcount == 523) begin
        // End of frame, reset counters
        hcount <= 0;
        vcount <= 0;
    end else if (hcount == 799) begin
        // End of line, reset hcount
        hcount <= 0;
        vcount <= vcount + 1;
    end else begin
        // Increment hcount
        hcount <= hcount + 1;
    end

    // Update sync and blanking signals
    hblank <= next_hblank;
    hsync <= hsyncon ? 0 : hsyncoff ? 1 : hsync;  // active low
    vblank <= next_vblank;
    vsync <= vsyncon ? 0 : vsyncoff ? 1 : vsync;  // active low
    blank <= next_vblank | (next_hblank & ~hreset);
end

endmodule