module karnaugh_map(
  input wire A, B, C, D, E,
  output reg F
);

always @(*) begin
  case ({A,B,C,D,E})
    5'b00000: F = 1;
    5'b00001: F = 0;
    5'b00011: F = 0;
    5'b00010: F = 0;
    5'b00110: F = 0;
    5'b00111: F = 1;
    5'b00101: F = 1;
    5'b00100: F = 0;
    5'b01100: F = 0;
    5'b01101: F = 1;
    5'b01111: F = 1;
    5'b01110: F = 1;
    5'b01010: F = 1;
    5'b01011: F = 1;
    5'b01001: F = 1;
    5'b01000: F = 0;
    5'b11000: F = 1;
    5'b11001: F = 0;
    5'b11011: F = 0;
    5'b11010: F = 0;
    5'b11110: F = 1;
    5'b11111: F = 1;
    5'b11101: F = 0;
    5'b11100: F = 0;
    5'b10100: F = 0;
    5'b10101: F = 0;
    5'b10111: F = 0;
    5'b10110: F = 0;
    5'b10010: F = 1;
    5'b10011: F = 1;
    5'b10001: F = 0;
    5'b10000: F = 0;
    default: F = 0;
  endcase
end

endmodule