module combinational_circuit (
    input A1,
    input A2,
    input A3,
    input B1,
    input B2,
    output X
);

    // Voltage supply signals
    supply1 VPWR;
    supply0 VGND;
    supply1 VPB ;
    supply0 VNB ;

    assign X = (A1 == 1'b1) ? B1 : ((A2 == 1'b1) && (A3 == 1'b0)) ? B2 : B1;

endmodule