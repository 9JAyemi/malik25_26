module StateUpdater(clk, enable, code, addr, state);

input clk, enable;
input [6:0] addr;
input [6:0] code;
output reg [3:0] state;

always @(posedge clk) begin
    if (enable) begin
        case (code)
            7'b0000000: state <= 4'b0000; // all 0s
            7'b1111111: state <= 4'b1111; // all 1s
            7'bxxxxxx1: state <= state ^ (1 << addr); // toggle
            7'bxxxxx1x: state <= state | (1 << addr); // set to 1
            7'bxxxx1xx: state <= state & ~(1 << addr); // set to 0
            7'bxxx1xxx: state <= state ^ (1 << addr); // invert
            7'bxx1xxxx: state <= {state[2:0], 1'b0}; // left shift
            7'bx1xxxxx: state <= {1'b0, state[3:1]}; // right shift
        endcase
    end
end

endmodule