module font_decoder(
    input wire [31:0] font_data_in,
    output reg [27:0] seg_out
);

    always @(*) begin
        case(font_data_in)
            4'b0000_0000_0000_0000_0000_0000_0000_0001: seg_out = {7'b0111111, 7'b0000110, 7'b1011011, 7'b1001111};
            4'b0000_0000_0000_0000_0000_0000_0000_0010: seg_out = {7'b0000110, 7'b0000110, 7'b1111101, 7'b0000111};
            4'b0000_0000_0000_0000_0000_0000_0000_0011: seg_out = {7'b1011011, 7'b0000110, 7'b1101101, 7'b1001111};
            4'b0000_0000_0000_0000_0000_0000_0000_0100: seg_out = {7'b1001110, 7'b1100110, 7'b0000110, 7'b0000111};
            4'b0000_0000_0000_0000_0000_0000_0000_0101: seg_out = {7'b1111101, 7'b1101101, 7'b0000110, 7'b1001111};
            4'b0000_0000_0000_0000_0000_0000_0000_0110: seg_out = {7'b1111111, 7'b1101101, 7'b0000110, 7'b1001111};
            4'b0000_0000_0000_0000_0000_0000_0000_0111: seg_out = {7'b0000111, 7'b0000110, 7'b1011011, 7'b0000111};
            4'b0000_0000_0000_0000_0000_0000_0000_1000: seg_out = {7'b1111111, 7'b1101111, 7'b0000110, 7'b1001111};
            4'b0000_0000_0000_0000_0000_0000_0000_1001: seg_out = {7'b1111101, 7'b1101101, 7'b0000110, 7'b1001111};
            default: seg_out = 28'b0;
        endcase
    end

endmodule