module Instruction_Mem(Instruction_out, PCAdress);
  output reg [15:0] Instruction_out;
  input  [15:0] PCAdress;
  
  always @(PCAdress)
  begin
    case (PCAdress)
 
		8'h0:  Instruction_out = 16'hc000; 8'h1:  Instruction_out = 16'ha802; 8'h2:  Instruction_out = 16'hc66b; 8'h3:  Instruction_out = 16'hec00; 8'h4:  Instruction_out = 16'hd119; 8'h5:  Instruction_out = 16'h6895; 8'h6:  Instruction_out = 16'h6805; 8'h7:  Instruction_out = 16'h696d; 8'h8:  Instruction_out = 16'h68aa; 8'h9:  Instruction_out = 16'h7168; 8'ha:  Instruction_out = 16'h6805; 8'hb:  Instruction_out = 16'h7168; 8'hc:  Instruction_out = 16'h6895; 8'hd:  Instruction_out = 16'h6368; 8'he:  Instruction_out = 16'h6802; 8'hf:  Instruction_out = 16'h6802; 8'h10:  Instruction_out = 16'ha818; 8'h11:  Instruction_out = 16'haa19; 8'h12:  Instruction_out = 16'had1a; 8'h13:  Instruction_out = 16'hf014; 8'h14:  Instruction_out = 16'ha003; 8'h15:  Instruction_out = 16'h4640; 8'h16:  Instruction_out = 16'h1901; 8'h17:  Instruction_out = 16'hb108; 8'h18:  Instruction_out = 16'h4640; 8'h19:  Instruction_out = 16'h1902; 8'h1a:  Instruction_out = 16'hb110; 8'h1b:  Instruction_out = 16'h4640; 8'h1c:  Instruction_out = 16'h1904; 8'h1d:  Instruction_out = 16'hb119; 8'h1e:  Instruction_out = 16'h9b80; 8'h1f:  Instruction_out = 16'hc000; 8'h20:  Instruction_out = 16'h5840; 8'h21:  Instruction_out = 16'h5888; 8'h22:  Instruction_out = 16'h58d0; 8'h23:  Instruction_out = 16'h5918; 8'h24:  Instruction_out = 16'h5960; 8'h25:  Instruction_out = 16'ha703; 8'h26:  Instruction_out = 16'h47f8; 8'h27:  Instruction_out = 16'h1f01; 8'h28:  Instruction_out = 16'hb7fd; 8'h29:  Instruction_out = 16'h9b80; 8'h2a:  Instruction_out = 16'hc000; 8'h2b:  Instruction_out = 16'h6400; 8'h2c:  Instruction_out = 16'h5840; 8'h2d:  Instruction_out = 16'h5888; 8'h2e:  Instruction_out = 16'h58d0; 8'h2f:  Instruction_out = 16'h5918; 8'h30:  Instruction_out = 16'h5960; 8'h31:  Instruction_out = 16'ha703; 8'h32:  Instruction_out = 16'h47f8; 8'h33:  Instruction_out = 16'h1f02; 8'h34:  Instruction_out = 16'hb7fd; 8'h35:  Instruction_out = 16'h9b80; 8'h36:  Instruction_out = 16'ha018; 8'h37:  Instruction_out = 16'ha219; 8'h38:  Instruction_out = 16'ha51a; 8'h39:  Instruction_out = 16'h5850; 8'h3a:  Instruction_out = 16'h2940; 8'h3b:  Instruction_out = 16'hf808; 8'h3c:  Instruction_out = 16'h6c4f; 8'h3d:  Instruction_out = 16'hf801; 8'h3e:  Instruction_out = 16'h4ccf; 8'h3f:  Instruction_out = 16'h6cdd; 8'h40:  Instruction_out = 16'h5900; 8'h41:  Instruction_out = 16'he800; 8'h42:  Instruction_out = 16'ha703; 8'h43:  Instruction_out = 16'h47f8; 8'h44:  Instruction_out = 16'h1f04; 8'h45:  Instruction_out = 16'hb7fd; 8'h46:  Instruction_out = 16'h9b80; 


		
	







      default: Instruction_out = 16'b0000000000000000;
    endcase
  end
endmodule 
