module adder32 ( 
    a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15,
    b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15,
    s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15,
    cout  );
  input  a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, 
b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15;
  output s0, s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13, s14, s15, cout;
  wire n50, n51, n53, n54, n55, n56, n57, n58, n60, n61, n62, n63, n64, n65,    n66, n67, n68, n69, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,    n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96,    n97, n98, n99, n100, n101, n102, n104, n105, n106, n107, n108, n109,    n110, n111, n112, n113, n115, n116, n117, n118, n119, n120, n121, n122,    n123, n124, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n148, n149,    n150, n151, n152, n153, n154, n155, n156, n157, n159, n160, n161, n162,    n163, n164, n165, n166, n167, n168, n170, n171, n172, n173, n174, n175,    n176, n177, n178, n179, n181, n182, n183, n184, n185, n186, n187, n188,    n189, n190, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,    n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n214, n215,   n216, n217;
  assign n50 = ~a0 & b0;
  assign n51 = a0 & ~b0;
  assign s0 = n50 | n51;
  assign n53 = a0 & b0;
  assign n54 = ~a1 & b1;
  assign n55 = a1 & ~b1;
  assign n56 = ~n54 & ~n55;
  assign n57 = n53 & n56;
  assign n58 = ~n53 & ~n56;
  assign s1 = n57 | n58;
  assign n60 = a1 & b1;
  assign n61 = a1 & n53;
  assign n62 = ~n60 & ~n61;
  assign n63 = b1 & n53;
  assign n64 = n62 & ~n63;
  assign n65 = ~a2 & b2;
  assign n66 = a2 & ~b2;
  assign n67 = ~n65 & ~n66;
  assign n68 = ~n64 & n67;
  assign n69 = n64 & ~n67;
  assign s2 = n68 | n69;
  assign n71 = a2 & b2;
  assign n72 = a2 & ~n64;
  assign n73 = ~n71 & ~n72;
  assign n74 = b2 & ~n64;
  assign n75 = n73 & ~n74;
  assign n76 = ~a3 & b3;
  assign n77 = a3 & ~b3;
  assign n78 = ~n76 & ~n77;
  assign n79 = ~n75 & n78;
  assign n80 = n75 & ~n78;
  assign s3 = n79 | n80;
  assign n82 = a3 & b3;
  assign n83 = a3 & ~n75;
  assign n84 = ~n82 & ~n83;
  assign n85 = b3 & ~n75;
  assign n86 = n84 & ~n85;
  assign n87 = ~a4 & b4;
  assign n88 = a4 & ~b4;
  assign n89 = ~n87 & ~n88;
  assign n90 = ~n86 & n89;
  assign n91 = n86 & ~n89;
  assign s4 = n90 | n91;
  assign n93 = a4 & b4;
  assign n94 = a4 & ~n86;
  assign n95 = ~n93 & ~n94;
  assign n96 = b4 & ~n86;
  assign n97 = n95 & ~n96;
  assign n98 = ~a5 & b5;
  assign n99 = a5 & ~b5;
  assign n100 = ~n98 & ~n99;
  assign n101 = ~n97 & n100;
  assign n102 = n97 & ~n100;
  assign s5 = n101 | n102;
  assign n104 = a5 & b5;
  assign n105 = a5 & ~n97;
  assign n106 = ~n104 & ~n105;
  assign n107 = b5 & ~n97;
  assign n108 = n106 & ~n107;
  assign n109 = ~a6 & b6;
  assign n110 = a6 & ~b6;
  assign n111 = ~n109 & ~n110;
  assign n112 = ~n108 & n111;
  assign n113 = n108 & ~n111;
  assign s6 = n112 | n113;
  assign n115 = a6 & b6;
  assign n116 = a6 & ~n108;
  assign n117 = ~n115 & ~n116;
  assign n118 = b6 & ~n108;
  assign n119 = n117 & ~n118;
  assign n120 = ~a7 & b7;
  assign n121 = a7 & ~b7;
  assign n122 = ~n120 & ~n121;
  assign n123 = ~n119 & n122;
  assign n124 = n119 & ~n122;
  assign s7 = n123 | n124;
  assign n126 = a7 & b7;
  assign n127 = a7 & ~n119;
  assign n128 = ~n126 & ~n127;
  assign n129 = b7 & ~n119;
  assign n130 = n128 & ~n129;
  assign n131 = ~a8 & b8;
  assign n132 = a8 & ~b8;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~n130 & n133;
  assign n135 = n130 & ~n133;
  assign s8 = n134 | n135;
  assign n137 = a8 & b8;
  assign n138 = a8 & ~n130;
  assign n139 = ~n137 & ~n138;
  assign n140 = b8 & ~n130;
  assign n141 = n139 & ~n140;
  assign n142 = ~a9 & b9;
  assign n143 = a9 & ~b9;
  assign n144 = ~n142 & ~n143;
  assign n145 = ~n141 & n144;
  assign n146 = n141 & ~n144;
  assign s9 = n145 | n146;
  assign n148 = a9 & b9;
  assign n149 = a9 & ~n141;
  assign n150 = ~n148 & ~n149;
  assign n151 = b9 & ~n141;
  assign n152 = n150 & ~n151;
  assign n153 = ~a10 & b10;
  assign n154 = a10 & ~b10;
  assign n155 = ~n153 & ~n154;
  assign n156 = ~n152 & n155;
  assign n157 = n152 & ~n155;
  assign s10 = n156 | n157;
  assign n159 = a10 & b10;
  assign n160 = a10 & ~n152;
  assign n161 = ~n159 & ~n160;
  assign n162 = b10 & ~n152;
  assign n163 = n161 & ~n162;
  assign n164 = ~a11 & b11;
  assign n165 = a11 & ~b11;
  assign n166 = ~n164 & ~n165;
  assign n167 = ~n163 & n166;
  assign n168 = n163 & ~n166;
  assign s11 = n167 | n168;
  assign n170 = a11 & b11;
  assign n171 = a11 & ~n163;
  assign n172 = ~n170 & ~n171;
  assign n173 = b11 & ~n163;
  assign n174 = n172 & ~n173;
  assign n175 = ~a12 & b12;
  assign n176 = a12 & ~b12;
  assign n177 = ~n175 & ~n176;
  assign n178 = ~n174 & n177;
  assign n179 = n174 & ~n177;
  assign s12 = n178 | n179;
  assign n181 = a12 & b12;
  assign n182 = a12 & ~n174;
  assign n183 = ~n181 & ~n182;
  assign n184 = b12 & ~n174;
  assign n185 = n183 & ~n184;
  assign n186 = ~a13 & b13;
  assign n187 = a13 & ~b13;
  assign n188 = ~n186 & ~n187;
  assign n189 = ~n185 & n188;
  assign n190 = n185 & ~n188;
  assign s13 = n189 | n190;
  assign n192 = a13 & b13;
  assign n193 = a13 & ~n185;
  assign n194 = ~n192 & ~n193;
  assign n195 = b13 & ~n185;
  assign n196 = n194 & ~n195;
  assign n197 = ~a14 & b14;
  assign n198 = a14 & ~b14;
  assign n199 = ~n197 & ~n198;
  assign n200 = ~n196 & n199;
  assign n201 = n196 & ~n199;
  assign s14 = n200 | n201;
  assign n203 = a14 & b14;
  assign n204 = a14 & ~n196;
  assign n205 = ~n203 & ~n204;
  assign n206 = b14 & ~n196;
  assign n207 = n205 & ~n206;
  assign n208 = ~a15 & b15;
  assign n209 = a15 & ~b15;
  assign n210 = ~n208 & ~n209;
  assign n211 = ~n207 & n210;
  assign n212 = n207 & ~n210;
  assign s15 = n211 | n212;
  assign n214 = a15 & b15;
  assign n215 = a15 & ~n207;
  assign n216 = ~n214 & ~n215;
  assign n217 = b15 & ~n207;
  assign cout = ~n216 | n217;
endmodule


