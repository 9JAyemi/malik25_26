module inverter (
    input A,
    output Y
);

    // Voltage supply signals
    supply1 VPWR;
    supply0 VGND;

    // Define internal signals
    wire A_valid;
    wire A_low;
    wire A_high;

    // Check if A is a valid logic level
    assign A_valid = (A == 0 || A == 1);

    // Check if A is low or high
    assign A_low = (A == 0);
    assign A_high = (A == 1);

    // Define the inverter logic
    assign Y = A_valid ? ~A : 1'bx;

endmodule