
module parity_generator (
    input [7:0] data_in,
    output reg parity_out
);

    always @(*) begin
        case (data_in)
            8'b00000001, 8'b00000011, 8'b00000101, 8'b00000111,
            8'b00001001, 8'b00001011, 8'b00001101, 8'b00001111,
            8'b00010001, 8'b00010011, 8'b00010101, 8'b00010111,
            8'b00011001, 8'b00011011, 8'b00011101, 8'b00011111,
            8'b00100001, 8'b00100011, 8'b00100101, 8'b00100111,
            8'b00101001, 8'b00101011, 8'b00101101, 8'b00101111,
            8'b00110001, 8'b00110011, 8'b00110101, 8'b00110111,
            8'b00111001, 8'b00111011, 8'b00111101, 8'b00111111,
            8'b01000001, 8'b01000011, 8'b01000101, 8'b01000111,
            8'b01001001, 8'b01001011, 8'b01001101, 8'b01001111,
            8'b01010001, 8'b01010011, 8'b01010101, 8'b01010111,
            8'b01011001, 8'b01011011, 8'b01011101, 8'b01011111,
            8'b01100001, 8'b01100011, 8'b01100101, 8'b01100111,
            8'b01101001, 8'b01101011, 8'b01101101, 8'b01101111,
            8'b01110001, 8'b01110011, 8'b01110101, 8'b01110111,
            8'b01111001, 8'b01111011, 8'b01111101, 8'b01111111,
            8'b10000001, 8'b10000011, 8'b10000101, 8'b10000111,
            8'b10001001, 8'b10001011, 8'b10001101, 8'b10001111,
            8'b10010001, 8'b10010011, 8'b10010101, 8'b10010111,
            8'b10011001, 8'b10011011, 8'b10011101, 8'b10011111,
            8'b10100001, 8'b10100011, 8'b10100101, 8'b10100111,
            8'b10101001, 8'b10101011, 8'b10101101, 8'b10101111,
            8'b10110001, 8'b10110011, 8'b10110101, 8'b10110111,
            8'b10111001, 8'b10111011, 8'b10111101, 8'b10111111,
            8'b11000001, 8'b11000011, 8'b11000101, 8'b11000111,
            8'b11001001, 8'b11001011, 8'b11001101, 8'b11001111,
            8'b11010001, 8'b11010011, 8'b11010101, 8'b11010111,
            8'b11011001, 8'b11011011, 8'b11011101, 8'b11011111,
            8'b11100001, 8'b11100011, 8'b11100101, 8'b11100111,
            8'b11101001, 8'b11101011, 8'b11101101, 8'b11101111,
            8'b11110001, 8'b11110011, 8'b11110101, 8'b11110111,
            8'b11111001, 8'b11111011, 8'b11111101, 8'b11111111:
                parity_out = 1;
            default:
                parity_out = 0;
        endcase
    end

endmodule

module parity_byte (
    input clk,
    input reset,
    input [7:0] a,
    input [7:0] b,
    input sel_b1,
    input sel_b2,
    output reg [8:0] out_byte
);

    reg [7:0] data_in;
    wire parity_out;

    // 2-to-1 mux to select between a and b
    always @(*) begin
        if (sel_b1 == 1 && sel_b2 == 0) begin
            data_in = a;
        end else if (sel_b1 == 0 && sel_b2 == 1) begin
            data_in = b;
        end else begin
            data_in = 8'b0;
        end
    end

    // Priority encoder to generate parity bit
    parity_generator parity (
        .data_in(data_in),
        .parity_out(parity_out)
    );

    // Multiplexer to combine parity bit and original 8 data bits
    always @(*) begin
        out_byte = {parity_out, data_in};
    end

endmodule
