module shift_register (
    in,
    shift,
    reset,
    clk,
    out
);

input [7:0] in;
input shift, reset, clk;
output [7:0] out;

reg [7:0] shift_reg;

always @ (posedge clk or posedge reset) begin
    if (reset) begin
        shift_reg <= 8'b0;
    end else if (shift) begin
        shift_reg <= {shift_reg[6:0], in};
    end
end

assign out = shift_reg;

endmodule