



module var6_multi(A, B, C, D, E, F, valid);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  
  input A;
  
  input B;
  
  input C;
  
  input D;
  
  input E;
  
  input F;
  
  wire [7:0] total_value;
  
  output valid;
  assign _43_ = C & D;
  assign _44_ = _43_ ^ A;
  assign _00_ = ~E;
  assign _01_ = ~(C | D);
  assign _02_ = ~(_01_ | _00_);
  assign _03_ = ~(_02_ & _44_);
  assign _04_ = ~(A ^ B);
  assign _05_ = ~(A & D);
  assign _06_ = _05_ & C;
  assign _07_ = _06_ ^ _04_;
  assign _08_ = _07_ | _00_;
  assign _09_ = _08_ & _03_;
  assign _10_ = ~D;
  assign _11_ = ~B;
  assign _12_ = A | _11_;
  assign _13_ = A & _11_;
  assign _14_ = ~((_13_ | C) & _12_);
  assign _15_ = _14_ & _10_;
  assign _16_ = ~(_14_ | _10_);
  assign _17_ = A & B;
  assign _18_ = ~(_17_ & C);
  assign _19_ = ~((_18_ & _16_) | _15_);
  assign _20_ = _19_ ^ _00_;
  assign _21_ = _20_ ^ _09_;
  assign _22_ = ~F;
  assign _23_ = _03_ & E;
  assign _24_ = _23_ ^ _07_;
  assign _25_ = E ? _43_ : _01_;
  assign _26_ = ~(_02_ | _44_);
  assign _27_ = _26_ & _25_;
  assign _28_ = ~((_27_ & _24_) | _22_);
  assign _29_ = _28_ | _21_;
  assign _30_ = _14_ | _10_;
  assign _31_ = A | B;
  assign _32_ = ~((_17_ | C) & _31_);
  assign _33_ = ~((_32_ & _30_) | (_43_ & A));
  assign _34_ = ~((_19_ & E) | _33_);
  assign _35_ = ~((_20_ | _09_) & _34_);
  assign _36_ = _26_ | _25_;
  assign _37_ = ~((_36_ | _24_) & _22_);
  assign _38_ = _37_ & _35_;
  assign _39_ = A | _10_;
  assign _40_ = _39_ | _22_;
  assign _41_ = E ? C : _11_;
  assign _42_ = _41_ | _40_;
  assign valid = ~((_38_ & _29_) | _42_);
  assign total_value[1:0] = { E, 1'b0 };
endmodule
