`define REGISTER_READ_OPERATION 1
`define REGISTER_WRITE_OPERATION 2


    module axi_slave_impl #
    (
        parameter integer NUMBER_OF_REGISTERS = 16,
        parameter integer C_S_AXI_DATA_WIDTH = 32,
        parameter integer C_S_AXI_ADDR_WIDTH = 10
    )
    (
        input wire [1:0] register_operation,      input wire [7 : 0] register_number,
		input wire [C_S_AXI_DATA_WIDTH -1 : 0] register_write,
		output reg [C_S_AXI_DATA_WIDTH -1 : 0] register_read,
        input wire S_AXI_ACLK,
        input wire S_AXI_ARESETN,
        input wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
        input wire [2 : 0] S_AXI_AWPROT,
        input wire  S_AXI_AWVALID,
        output wire  S_AXI_AWREADY,
        input wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_WDATA,
        input wire [(C_S_AXI_DATA_WIDTH/8)-1 : 0] S_AXI_WSTRB,
        input wire  S_AXI_WVALID,
        output wire  S_AXI_WREADY,
        output wire [1 : 0] S_AXI_BRESP,
        output wire  S_AXI_BVALID,
        input wire  S_AXI_BREADY,
        input wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
        input wire [2 : 0] S_AXI_ARPROT,
        input wire  S_AXI_ARVALID,
        output wire  S_AXI_ARREADY,
        output wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_RDATA,
        output wire [1 : 0] S_AXI_RRESP,
        output wire  S_AXI_RVALID,
        input wire  S_AXI_RREADY
    );

     reg [C_S_AXI_ADDR_WIDTH-1 : 0] axi_awaddr;
    reg axi_awready;
    reg axi_wready;
     reg [1 : 0] axi_bresp;
    reg axi_bvalid;
     reg [C_S_AXI_ADDR_WIDTH-1 : 0] axi_araddr;
    reg axi_arready;
    reg [C_S_AXI_DATA_WIDTH-1 : 0] axi_rdata;
     reg [1 : 0] axi_rresp;
    reg axi_rvalid;

    localparam integer ADDR_LSB = (C_S_AXI_DATA_WIDTH/32) + 1;
    localparam integer OPT_MEM_ADDR_BITS =  C_S_AXI_ADDR_WIDTH - ADDR_LSB - 1;
    reg register_operation_done;
    reg [C_S_AXI_DATA_WIDTH-1:0] registers[NUMBER_OF_REGISTERS - 1 : 0];
    wire slv_reg_rden;
    wire slv_reg_wren;
    reg [C_S_AXI_DATA_WIDTH-1:0] reg_data_out;
    integer byte_index;
    integer register_index;
    assign S_AXI_AWREADY = axi_awready;
    assign S_AXI_WREADY = axi_wready;
    assign S_AXI_BRESP = axi_bresp;
    assign S_AXI_BVALID = axi_bvalid;
    assign S_AXI_ARREADY = axi_arready;
    assign S_AXI_RDATA = axi_rdata;
    assign S_AXI_RRESP = axi_rresp;
    assign S_AXI_RVALID = axi_rvalid;
    
    always @(posedge S_AXI_ACLK)
    begin
        if (S_AXI_ARESETN == 1'b0)
        begin
            axi_awready <= 1'b0;
        end 
        else
        begin    
            if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID)
            begin
                axi_awready <= 1'b1;
            end
            else           
            begin
                axi_awready <= 1'b0;
            end
        end 
    end       

    always @(posedge S_AXI_ACLK)
    begin
        if (S_AXI_ARESETN == 1'b0)
        begin
            axi_awaddr <= 0;
        end 
        else
        begin    
            if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID)
            begin
                axi_awaddr <= S_AXI_AWADDR;
            end
        end 
    end       

    always @(posedge S_AXI_ACLK)
    begin
        if (S_AXI_ARESETN == 1'b0)
        begin
            axi_wready <= 1'b0;
        end 
        else
        begin    
            if (~axi_wready && S_AXI_WVALID && S_AXI_AWVALID)
            begin
                axi_wready <= 1'b1;
            end
            else
            begin
                axi_wready <= 1'b0;
            end
        end 
    end       

    assign slv_reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;

    always @(posedge S_AXI_ACLK)
    begin
        if (S_AXI_ARESETN == 1'b0)
        begin
            for (register_index = 0; register_index < NUMBER_OF_REGISTERS; register_index = register_index + 1)
                registers[register_index] <= 0;
        end 
        else 
        if (slv_reg_wren)
        begin
             for (byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH / 8) -1; byte_index = byte_index + 1)
             begin
                 if (S_AXI_WSTRB[byte_index] == 1) 
                     registers[axi_awaddr[ADDR_LSB + OPT_MEM_ADDR_BITS : ADDR_LSB]][(byte_index * 8) +: 8] <= S_AXI_WDATA[(byte_index * 8) +: 8];
             end
        end
		else
		begin
		    if(register_operation == `REGISTER_WRITE_OPERATION && register_number > 0)
		    begin
		        registers[register_number - 1] <= register_write;
		    end
		end
    end    

    always @(posedge S_AXI_ACLK)
    begin
        if (S_AXI_ARESETN == 1'b0)
        begin
            axi_bvalid  <= 0;
            axi_bresp   <= 2'b0;
        end 
        else
        begin    
            if (axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID)
            begin
                axi_bvalid <= 1'b1;
                axi_bresp  <= 2'b0; end                   else
            begin
                if (S_AXI_BREADY && axi_bvalid) 
				begin
                axi_bvalid <= 1'b0; 
                end  
            end
        end
    end   

    always @(posedge S_AXI_ACLK)
    begin
        if (S_AXI_ARESETN == 1'b0)
        begin
            axi_arready <= 1'b0;
            axi_araddr  <= 32'b0;
        end 
        else
        begin    
            if (~axi_arready && S_AXI_ARVALID)
            begin
                axi_arready <= 1'b1;
                axi_araddr  <= S_AXI_ARADDR;
            end
            else
            begin
                axi_arready <= 1'b0;
            end
        end 
    end       

    always @(posedge S_AXI_ACLK)
    begin
        if ( S_AXI_ARESETN == 1'b0 )
        begin
            axi_rvalid <= 0;
            axi_rresp  <= 0;
        end 
        else
        begin    
            if (axi_arready && S_AXI_ARVALID && ~axi_rvalid)
            begin
                axi_rvalid <= 1'b1;
                axi_rresp  <= 2'b0; end   
            else if (axi_rvalid && S_AXI_RREADY)
            begin
                axi_rvalid <= 1'b0;
            end                
        end
    end    

    assign slv_reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;
    always @(*)
    begin
        if(axi_araddr[ADDR_LSB + OPT_MEM_ADDR_BITS : ADDR_LSB] < NUMBER_OF_REGISTERS)
           reg_data_out <= registers[axi_araddr[ADDR_LSB + OPT_MEM_ADDR_BITS : ADDR_LSB]];
        else reg_data_out <= 0;
    end

    always @(posedge S_AXI_ACLK)
    begin
        if (S_AXI_ARESETN == 1'b0)
        begin
            axi_rdata  <= 0;
        end 
        else
        begin    
            if (slv_reg_rden)
            begin
                axi_rdata <= reg_data_out;     end   
            else
            begin
                if(register_operation == `REGISTER_READ_OPERATION)
                begin
                    register_read <= registers[register_number - 1];
                    end
            end
        end
    end    

    endmodule
