module priority_encoder (
    input [3:0] I,
    output [15:0] O
);

    assign O = (I == 4'h0) ? 16'b0000000000000001 :
               (I == 4'h1) ? 16'b0000000000000010 :
               (I == 4'h2) ? 16'b0000000000000100 :
               (I == 4'h3) ? 16'b0000000000001000 :
               (I == 4'h4) ? 16'b0000000000010000 :
               (I == 4'h5) ? 16'b0000000000100000 :
               (I == 4'h6) ? 16'b0000000001000000 :
               (I == 4'h7) ? 16'b0000000010000000 :
               (I == 4'h8) ? 16'b0000000100000000 :
               (I == 4'h9) ? 16'b0000001000000000 :
               (I == 4'ha) ? 16'b0000010000000000 :
               (I == 4'hb) ? 16'b0000100000000000 :
               (I == 4'hc) ? 16'b0001000000000000 :
               (I == 4'hd) ? 16'b0010000000000000 :
               (I == 4'he) ? 16'b0100000000000000 :
                             16'b1000000000000000 ;

endmodule